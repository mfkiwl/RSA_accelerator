../lab3-qsys/VGA_LED_Emulator.sv