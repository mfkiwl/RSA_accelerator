../lab3-qsys/VGA_LED.sv