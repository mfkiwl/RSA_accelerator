/* verilator lint_off UNUSED */
module incrementA(input logic reset, input logic clk);
endmodule
