../lab3-qsys/RSA_BOX.sv